/*
Testbench for the General Controller FSM
*/
